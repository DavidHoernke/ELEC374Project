library verilog;
use verilog.vl_types.all;
entity registerTB is
end registerTB;
